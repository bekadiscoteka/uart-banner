`include "uart/uart.v"
`include "bcd2sseg_active_low.v"
`include "signal_decoder.v"
`include "serial2parallel.v"
`include "bcd_shift_register.v"
module top(
	output [7:0]	sseg5,
					sseg4,
					sseg3,
					sseg2,
					sseg1,
					sseg0,
	output	baund_rate_ready, //indicates baund is detected 
			banner_write, //indicates banner is being written
			tx,
	input clk, reset, rx
);				
	wire	rx_empty, read,
			write_banner,
			start,
			pause,
			left,
			right,
			s2p_done_tick;

	wire [7:0] ascii;
	wire [(4*6)-1:0] parallel_data, bcd_set;

	uart uart_inst(
		.clk(clk),
		.reset(reset),
		.rx(rx),
		.tx(tx),
		.data_in(),
		.data_out(ascii),
		.rx_empty(rx_empty), // rx fifo empty
		.ready(baund_rate_ready),
		.rd_data(read)
	);		

	assign read = ~rx_empty;

	signal_decoder dcode(
		.ascii(ascii),
		.write_banner(write_banner),
		.start(start),
		.pause(pause),
		.left(left),
		.right(right)
	);

	serial2parallel s2p(
		.clk(clk),
		.reset(reset),
		.start(write_banner),
		.new_in_data(!rx_empty),
		.done_tick(s2p_done_tick),
		.data_out(parallel_data),
		.data_in(ascii-48),
		.write_mode(banner_write)
	);

	bcd_shift_register sr(
		.clk(clk),
		.reset(reset),
		.set_left(left),
		.set_right(right),
		.start(start),
		.write(s2p_done_tick),
		.pause(pause),
		.data_in(parallel_data),
		.data_out(bcd_set)
	);

	bcd2sseg_active_low b2ssg(
		.bcd5(bcd_set[(4*6)-1:(4*6)-4]),
		.bcd4(bcd_set[(4*5)-1:(4*5)-4]),	
		.bcd3(bcd_set[(4*4)-1:(4*4)-4]),
		.bcd2(bcd_set[(4*3)-1:(4*3)-4]),
		.bcd1(bcd_set[(4*2)-1:(4*2)-4]),
		.bcd0(bcd_set[(4*1)-1:(4*1)-4]),
		.sseg5(sseg5[6:0]),
		.sseg4(sseg4[6:0]),
		.sseg3(sseg3[6:0]),
		.sseg2(sseg2[6:0]),
		.sseg1(sseg1[6:0]),
		.sseg0(sseg0[6:0])
	);	

	assign {sseg5[7], sseg4[7], sseg3[7], sseg2[7], sseg1[7], sseg0[7]} = ~6'b0;
	
endmodule
