Vim�UnDo� U��4�Z���e��5�v�f1��K����ce��u      	parameter DIVIDER=49_999      
                       h
G;    _�                            ����                                                                                                                                                                                                                                                                                                                                                             h�~     �                	input [25:0] divider5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             h�     �               module clk_div_26bit(5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             h�     �               	�             5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             h�     �               	parameter DIVIDER,5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             h�    �               	parameter DIVIDER5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             h�    �               $		else if (counter == divider) begin5�_�                    	       ����                                                                                                                                                                                                                                                                                                                                                             h��   	 �      
         	input clk, reset,5�_�                        
    ����                                                                                                                                                                                                                                                                                                                                                             h
G:    �               	parameter DIVIDER=49_9995��