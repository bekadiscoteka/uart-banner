Vim�UnDo� O��L�4q�1���8�dd&��`�EZb���    3                 �       �   �   �    h��   , _�                             ����                                                                                                                                                                                                                                                                                                                                                             h��     �                   5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             h��     �               	�             5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             h��     �               	module 5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             h�     �               		�             5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             h�     �               	module serial2parallel(5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             h�    �               		�             5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             h�J     �         	      			output 5�_�      	                     ����                                                                                                                                                                                                                                                                                                                                                             h�Y     �         	      		output [SERIAL_W-1:0] data 5�_�      
           	          ����                                                                                                                                                                                                                                                                                                                                                             h�`     �         	      (		output [SERIAL_W*PARALLEL_N-1:0] data 5�_�   	              
      
    ����                                                                                                                                                                                                                                                                                                                                                             h�c     �         	      )		output [SERIAL_W*PARALLEL_N)-1:0] data 5�_�   
                    *    ����                                                                                                                                                                                                                                                                                                                                                             h�{     �      	   	      *		output [(SERIAL_W*PARALLEL_N)-1:0] data 5�_�                       	    ����                                                                                                                                                                                                                                                                                                                                         	       v       h��     �      	   
      		input [PARALLEL_N-1:0]5�_�                       	    ����                                                                                                                                                                                                                                                                                                                                         	       v       h��     �      	   
      		input [-1:0]5�_�                           ����                                                                                                                                                                                                                                                                                                                                         	       v       h��     �      
   
      		input [SERIAL_W-1:0]5�_�                           ����                                                                                                                                                                                                                                                                                                                                         	       v       h��     �   
              `endif5�_�                    	       ����                                                                                                                                                                                                                                                                                                                                         	       v       h��     �               		input clk, reset, 5�_�                    
        ����                                                                                                                                                                                                                                                                                                                                         	       v       h��     �   	   
           5�_�                    	   "    ����                                                                                                                                                                                                                                                                                                                                         	       v       h��     �      
         "		input clk, reset, write_tick_in,5�_�                            ����                                                                                                                                                                                                                                                                                                                                         	       v       h��    �      	         		�      	       5�_�                           ����                                                                                                                                                                                                                                                                                                                            	          	   	       v       h��     �               		�             5�_�                           ����                                                                                                                                                                                                                                                                                                                            	          	   	       v       h��     �             5�_�                            ����                                                                                                                                                                                                                                                                                                                            	          	   	       v       h��     �                5�_�                           ����                                                                                                                                                                                                                                                                                                                            	          	   	       v       h�     �               			�             5�_�                           ����                                                                                                                                                                                                                                                                                                                            	          	   	       v       h�	     �               				�             5�_�                           ����                                                                                                                                                                                                                                                                                                                            	          	   	       v       h�(    �               		�             5�_�                       
    ����                                                                                                                                                                                                                                                                                                                            	          	   	       v       h�K     �               					START;5�_�                           ����                                                                                                                                                                                                                                                                                                                            	          	   	       v       h�U     �               				5�_�                           ����                                                                                                                                                                                                                                                                                                                                                v       h�l     �               					CONVERT;5�_�                           ����                                                                                                                                                                                                                                                                                                                                                v       h�m     �               					;5�_�                           ����                                                                                                                                                                                                                                                                                                                                                v       h�o    �               					5�_�                            ����                                                                                                                                                                                                                                                                                                                                                v       h�{     �               				state <= 0;5�_�      !                      ����                                                                                                                                                                                                                                                                                                                                                v       h�~     �               			�             5�_�       $           !          ����                                                                                                                                                                                                                                                                                                                                                v       h��     �             5�_�   !   %   "       $           ����                                                                                                                                                                                                                                                                                                                                                v       h��     �                 5�_�   $   &           %          ����                                                                                                                                                                                                                                                                                                                                                v       h��     �               				�             5�_�   %   '           &      
    ����                                                                                                                                                                                                                                                                                                                                                v       h��     �               					�             5�_�   &   (           '          ����                                                                                                                                                                                                                                                                                                                                                v       h��     �               				�             5�_�   '   )           (      
    ����                                                                                                                                                                                                                                                                                                                                                v       h��    �               					IDLE: 5�_�   (   *           )      ,    ����                                                                                                                                                                                                                                                                                                                                                v       h��     �               					�             5�_�   )   +           *          ����                                                                                                                                                                                                                                                                                                                                                v       h��     �               						�             5�_�   *   ,           +   
   !    ����                                                                                                                                                                                                                                                                                                                                                v       h��    �   	            !		input clk, reset, write_tick_in5�_�   +   -           ,      
    ����                                                                                                                                                                                                                                                                                                                                                v       h��     �               
						if (5�_�   ,   .           -   
   #    ����                                                                                                                                                                                                                                                                                                                                                v       h��     �   	            3		input clk, reset, write_tick_in, special_ctrlwire5�_�   -   /           .          ����                                                                                                                                                                                                                                                                                                                                                v       h��     �   
             			  special_ctrlwire5�_�   .   0           /   
   "    ����                                                                                                                                                                                                                                                                                                                                                v       h��     �   	             #		input clk, reset, write_tick_in, 5�_�   /   1           0   
       ����                                                                                                                                                                                                                                                                                                                                                v       h��     �   	             $		input clk, reset, write_tick_in,  5�_�   0   2           1          ����                                                                                                                                                                                                                                                                                                                                                v       h��     �   
      !      			  write_tick_in,  5�_�   1   3           2          ����                                                                                                                                                                                                                                                                                                                                                v       h�     �         !      <			  special_ctrlwire // should be 1, at state of convertion5�_�   2   4           3          ����                                                                                                                                                                                                                                                                                                                                                v       h�      �         !      7			  new_data_in // should be 1, at state of convertion5�_�   3   5           4      	    ����                                                                                                                                                                                                                                                                                                                                                v       h�&     �         !      4			  new_data // should be 1, at state of convertion5�_�   4   6           5          ����                                                                                                                                                                                                                                                                                                                                                v       h�)     �   
      !      			  write_tick_in,  5�_�   5   7           6          ����                                                                                                                                                                                                                                                                                                                                                v       h�8     �   
      !      		write_tick_in,  //indicates 5�_�   6   8           7          ����                                                                                                                                                                                                                                                                                                                                                v       h�C     �   
      !      (		write_tick_in,  //indicates start of  5�_�   7   9           8          ����                                                                                                                                                                                                                                                                                                                                                v       h�G     �   
      !      +			  write_tick_in,  //indicates start of  5�_�   8   :           9          ����                                                                                                                                                                                                                                                                                                                                                v       h�H     �   
      !      			  ,  //indicates start of  5�_�   9   ;           :      #    ����                                                                                                                                                                                                                                                                                                                                                v       h�J     �   
      !      #			  start,  //indicates start of  5�_�   :   <           ;      7    ����                                                                                                                                                                                                                                                                                                                                                v       h�O     �         !      7			  new_in_data // should be 1, at state of convertion5�_�   ;   =           <          ����                                                                                                                                                                                                                                                                                                                                                v       h�_    �         !      1			  new_in_data // when there is new input data 5�_�   <   >           =      $    ����                                                                                                                                                                                                                                                                                                                                                v       h�e   	 �         !      3			  new_in_data // 1 when there is new input data 5�_�   =   ?           >          ����                                                                                                                                                                                                                                                                                                                                                v       h�y     �                						if (special_ctrlWire5�_�   >   @           ?          ����                                                                                                                                                                                                                                                                                                                                                v       h�z     �         !      						�              5�_�   ?   A           @          ����                                                                                                                                                                                                                                                                                                                                                v       h��     �         #      							�         "    5�_�   @   B           A          ����                                                                                                                                                                                                                                                                                                                                                v   *    h��     �         #      .					IDLE: if (write_tick_in) state <= START; 5�_�   A   C           B          ����                                                                                                                                                                                                                                                                                                                                                v   *    h��     �         #      !					IDLE: if () state <= START; 5�_�   B   D           C          ����                                                                                                                                                                                                                                                                                                                                                v   *    h��     �                							5�_�   C   E           D          ����                                                                                                                                                                                                                                                                                                                                                v   *    h��     �         #      							�         "    5�_�   D   F           E          ����                                                                                                                                                                                                                                                                                                                                                v   *    h��     �         #      							data_out <= {}5�_�   E   G           F           ����                                                                                                                                                                                                                                                                                                                                                v   *    h��     �      
           		input [SERIAL_W-1:0] data_in, �                .		output [(SERIAL_W*PARALLEL_N)-1:0] data_out,�                		parameter	SERIAL_W,5�_�   F   H           G           ����                                                                                                                                                                                                                                                                                                                                                v   *    h�    
 �                '		output [(W*PARALLEL_N)-1:0] data_out,�                					PARALLEL_N5�_�   G   I           H          ����                                                                                                                                                                                                                                                                                                                                                v   *    h�
     �         #      							data_out <= {}5�_�   H   J           I          ����                                                                                                                                                                                                                                                                                                                                                v   *    h�#     �         #      							data_out <= {W*N)}5�_�   I   K           J          ����                                                                                                                                                                                                                                                                                                                                                v   *    h�%     �         #      							data_out <= {(W*N)}5�_�   J   L           K          ����                                                                                                                                                                                                                                                                                                                                                v   *    h�;     �         #      							data_out <= {(W*N)-W)}5�_�   K   M           L          ����                                                                                                                                                                                                                                                                                                                                                v   *    h�=     �         #      							data_out <= {((W*N)-W)}5�_�   L   N           M          ����                                                                                                                                                                                                                                                                                                                                                v   *    h�?     �         #       							data_out <= {((W*N)-W){}}5�_�   M   O           N          ����                                                                                                                                                                                                                                                                                                                                                v   (    h�p     �         #       							data_out <= {((W*N)-W){}}5�_�   N   P           O          ����                                                                                                                                                                                                                                                                                                                                                v   (    h�r     �         #      							data_out <= 5�_�   O   Q           P          ����                                                                                                                                                                                                                                                                                                                                                v   (    h��     �         #      							data_out[W-1:0] <= 5�_�   P   R           Q          ����                                                                                                                                                                                                                                                                                                                                                v   (    h��    �         $      "							data_out[W-1:0] <= data_in;5�_�   Q   S           R           ����                                                                                                                                                                                                                                                                                                                                                v   (    h��     �         $       5�_�   R   T           S          ����                                                                                                                                                                                                                                                                                                                                                v   (    h��     �                				5�_�   S   U           T          ����                                                                                                                                                                                                                                                                                                                                                v   (    h��    �         $      							�         #    5�_�   T   V           U           ����                                                                                                                                                                                                                                                                                                                                                v   (    h��    �         %      							�         $    5�_�   U   W           V          ����                                                                                                                                                                                                                                                                                                                                                v   (    h�     �         &      							�         %    5�_�   V   X           W          ����                                                                                                                                                                                                                                                                                                                                                v   (    h�U     �         &      							if (counter == N-1)5�_�   W   Y           X      	    ����                                                                                                                                                                                                                                                                                                                                                v   (    h�X    �          (      								�         '    5�_�   X   Z           Y       	    ����                                                                                                                                                                                                                                                                                                                            !          !          v   (    h��     �       "   *    5�_�   Y   [           Z   "       ����                                                                                                                                                                                                                                                                                                                            "          $          v   2    h��     �   !   %   +      !							data_out[W-1:0] = data_in;   !							data_out <= data_out << W;   							counter <= counter + 1;5�_�   Z   \           [   !        ����                                                                                                                                                                                                                                                                                                                            "          $          v   2    h��     �       !           5�_�   [   ]           \       	    ����                                                                                                                                                                                                                                                                                                                            !          #          v   2    h��     �       "   +      							�       "   *    5�_�   \   ^           ]   $       ����                                                                                                                                                                                                                                                                                                                            "          $          v   2    h��    �   $   &   ,      								�   $   &   +    5�_�   ]   _           ^          ����                                                                                                                                                                                                                                                                                                                            "          $          v   2    h��    �          -      #								data_out[W-1:0] <= data_in;    �      !   -      								�      !   ,    5�_�   ^   `           _      
    ����                                                                                                                                                                                                                                                                                                                            "          $          v   2    h��     �         ,      &					IDLE: if (start) state <= START; 5�_�   _   a           `          ����                                                                                                                                                                                                                                                                                                                            #          %          v   2    h��     �         .      						�         -    5�_�   `   b           a          ����                                                                                                                                                                                                                                                                                                                            $          &          v   2    h��    �         /      						�         .    5�_�   a   c           b      
    ����                                                                                                                                                                                                                                                                                                                            '          )          v   2    h�     �         2      		�         1    5�_�   b   d           c          ����                                                                                                                                                                                                                                                                                                                            )          +          v   2    h�    �         3      		reg [N-1:0] 5�_�   c   e           d          ����                                                                                                                                                                                                                                                                                                                            *          ,          v   2    h�#    �         4    5�_�   d   f           e      
    ����                                                                                                                                                                                                                                                                                                                            +          -          v   2    h�'     �         5      					START;5�_�   e   g           f          ����                                                                                                                                                                                                                                                                                                                            +          -          v   2    h�)    �         5      		localparam	IDLE,5�_�   f   h           g          ����                                                                                                                                                                                                                                                                                                                            +          -          v   2    h�l     �      	   5      		output done_tick,5�_�   g   i           h          ����                                                                                                                                                                                                                                                                                                                            +          -          v   2    h�p    �         5      		output [(W*N)-1:0] data_out,5�_�   h   j           i          ����                                                                                                                                                                                                                                                                                                                            +          -          v   2    h��     �         5      		parameter	W,5�_�   i   k           j          ����                                                                                                                                                                                                                                                                                                                            +          -          v   2    h��    �         5      					N5�_�   j   l           k   +       ����                                                                                                                                                                                                                                                                                                                            5                     v        h�~     �   *   +          "								data_out[W-1:0] = data_in;5�_�   k   m           l   +       ����                                                                                                                                                                                                                                                                                                                            4                     v        h��     �   *   ,   4      "								data_out <= data_out << W;5�_�   l   n           m   +   "    ����                                                                                                                                                                                                                                                                                                                            4                     v        h��     �   *   ,   4      #								data_out <= (data_out << W;5�_�   m   o           n   +       ����                                                                                                                                                                                                                                                                                                                            4                     v        h��     �   *   ,   4      %								data_out <= (data_out << W) ;5�_�   n   p           o   +   #    ����                                                                                                                                                                                                                                                                                                                            4                     v        h��     �   *   ,   4      %								data_out <= (data_out << W) ;5�_�   o   q           p   +   $    ����                                                                                                                                                                                                                                                                                                                            4                     v        h��   ! �   *   ,   4      %								data_out <= (data_out << W) ;5�_�   p   s           q   $       ����                                                                                                                                                                                                                                                                                                                            +   -       +          v        h�     �   $   &   4    5�_�   q   t   r       s   %        ����                                                                                                                                                                                                                                                                                                                            ,   -       ,          v        h�     �   $   &   5       5�_�   s   u           t   %       ����                                                                                                                                                                                                                                                                                                                            ,   -       ,          v        h�     �   $   &   5      								�   %   &   5    5�_�   t   v           u   %       ����                                                                                                                                                                                                                                                                                                                            ,   -       ,          v        h�#   " �   $   &   5      .								data_out <= (data_out << W) | data_in;5�_�   u   w           v   ,       ����                                                                                                                                                                                                                                                                                                                            ,   -       ,          v        h�&     �   +   ,          .								data_out <= (data_out << W) | data_in;5�_�   v   x           w   -       ����                                                                                                                                                                                                                                                                                                                            ,   -       ,          v        h�,     �   ,   -          
							end5�_�   w   y           x   ,       ����                                                                                                                                                                                                                                                                                                                            ,   -       ,          v        h�-   # �   *   ,   3      							else begin   counter <= counter + 1;�   +   -   3      								counter <= counter + 1;5�_�   x   z           y   )       ����                                                                                                                                                                                                                                                                                                                            +   >       +          v        h�3   & �   (   )          #								data_out[W-1:0] <= data_in;5�_�   y   {           z          ����                                                                                                                                                                                                                                                                                                                            *   >       *          v        h�o     �         1      5			  new_in_data // 1 when there is a new input data 5�_�   z   |           {          ����                                                                                                                                                                                                                                                                                                                            *   >       *          v        h��   ' �         1      		parameter	W=8,5�_�   {   }           |   !       ����                                                                                                                                                                                                                                                                                                                            *   >       *          v        h��   ) �       !          						data_out <= 0;5�_�   |   ~           }          ����                                                                                                                                                                                                                                                                                                                            )   >       )          v        h��   * �      
   1      		�      
   0    5�_�   }              ~   	   	    ����                                                                                                                                                                                                                                                                                                                            	          	   	       v       h��     �      
   1      		output begin_written,5�_�   ~   �              	   	    ����                                                                                                                                                                                                                                                                                                                            	          	   	       v       h��   + �      
   1      
		output ,5�_�                  �          ����                                                                                                                                                                                                                                                                                                                            	          	   	       v       h��   , �         2      		�         1    5�_�   q           s   r   %        ����                                                                                                                                                                                                                                                                                                                            ,   -       ,          v        h�     �   %   &   5    �   $   &   5      &data_out <= (data_out << W) | data_in;5�_�   !   #       $   "           ����                                                                                                                                                                                                                                                                                                                                                v       h��     �               				case (state) begin   				end5�_�   "               #          ����                                                                                                                                                                                                                                                                                                                                                v       h��     �                5��